
context common_ctx is -- To be compiled in common_lib

    library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;

    use common_lib.logger_pkg.all;

end context;
